`define DATA_WIDTH 16

typedef enum {read, write} wr_rd_type ;
//typedef uvm_reg_predictor#(apb_transaction)  apb_predictor;   //map apb tx to register in model


