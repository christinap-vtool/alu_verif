
`timescale 1ns/100ps
`include "uvm_macros.svh"
`include "alu_interface.sv"
`include "alu_pkg.sv"
`include "alu_test_pkg.sv"
`include "top_tb.sv"

