`define DATA_WIDTH 16
`define DATA_SIZE 16
`define MUL_DATA_SIZE 8
`define FIFO_IN_DEPTH 4
`define FIFO_OUT_DEPTH 4
`define APB_BUS_SIZE 32
`define REG_NUMBER 5

typedef enum {read, write} wr_rd_type ;


