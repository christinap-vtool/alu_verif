`define DATA_WIDTH 16
`define DATA_SIZE 16           //todo maybe should be found only in the defines
`define MUL_DATA_SIZE 8
`define FIFO_IN_DEPTH 4
`define FIFO_OUT_DEPTH 4

typedef enum {read, write} wr_rd_type ;


